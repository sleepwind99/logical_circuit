`timescale 1ns/1ps

module SAM();
  reg clk;

// TODO: you may alter the type of registers to wire (e.g. reg RW -> wire RW) if necessary
  reg [15:0] PC;
  reg [15:0] AC, MAR, MBR, IR;
  reg [15:0] ABUS, RBUS, MBUS;
  reg [15:0] ADDRESS_BUS, DATA_BUS;
  reg RW, REQUEST;
  wire WAIT;

  reg [15:0] ALU_A, ALU_B;
  reg ALU_ADD, ALU_PASS_B;
  reg [15:0] ALU_RESULT;

  wire [21:0] b;
  controller my_controller(clk, WAIT, IR[15], AC[15], IR[14], b);

  wire [15:0] data_bus_t;
  always @ ( RW ) if (RW) DATA_BUS = data_bus_t;
  Memory my_memory(ADDRESS_BUS, REQUEST, RW, WAIT, DATA_BUS, data_bus_t);

  // initial settings
  // TODO : add any initialization process if required (not necessary)
  initial begin
    clk = 0;
    AC = 0;
    IR = 0;
    ADDRESS_BUS = 0;
  end
  always begin
    clk = ~clk; #1;
  end

  // ALU implementation
  always @ (ALU_ADD or ALU_PASS_B or ALU_A or ALU_B )begin
    if (ALU_ADD) ALU_RESULT = ALU_A + ALU_B;
    else if (ALU_PASS_B) ALU_RESULT = ALU_B;
  end

  always @ ( negedge clk ) begin
  // TODO: refer to lecture note, page 46
   if (b[21]) ABUS = PC; //b21
   if (b[20]) ABUS = IR; //b20
   if (b[19]) ABUS = MBR; //b19
   if (b[7]) MBUS = MBR; //b7
   if (b[16]) ALU_B = MBUS; //b16
   if (b[14]) begin //b14
    ALU_PASS_B = 1;
    ALU_RESULT = ALU_B;
   end
   else ALU_PASS_B = 0;
   if (b[0]) RBUS = ALU_RESULT; //b0
   if (b[18]) AC = RBUS; //b18
   if (b[17]) ALU_A = AC; //b17
   if (b[15]) begin //b15
    ALU_ADD = 1; 
   end
 	 else ALU_ADD = 0;
   if (b[13]) ADDRESS_BUS = MAR; //b13
   if (b[12]) DATA_BUS = MBR; //b12
   if (b[11]) IR = ABUS; //b11
   if (b[10]) MAR = ABUS; //b10
   if (b[9]) MBR = DATA_BUS; //b9
   if (b[8]) MBR = RBUS; //b8
   if (b[6]) PC = 0; //b6
   if (b[5]) PC = PC+2; //b5
   if (b[4]) PC = ABUS; //b4
   if (b[3]) begin //b3
    RW = 1;
   end
   else RW = 0;
   if (b[2]) begin //b2
    REQUEST = 1; 
   end
   else REQUEST = 0;
   if (b[1]) RBUS = AC; //b1
  end
 
  //always @ (b or PC or IR or MBR) begin
//    if (b[19]) ABUS = MBR; //b19
//    if (b[18]) AC = RBUS; //b18
//    if (b[17]) ALU_A = AC; //b17
//    if (b[16]) ALU_B = MBUS; //b16
//    if (b[15]) begin //b15
//    ALU_ADD = 1; 
//    end
//   	else ALU_ADD = 0;
//    if (b[14]) begin //b14
//    ALU_PASS_B = 1; 
//    end
//    else ALU_PASS_B = 0; 
//    if (b[11]) IR = ABUS; //b11
//    if (b[10]) MAR = ABUS; //b10
//    if (b[7]) MBUS = MBR; //b7
//    if (b[6]) PC = 0; //b6
//    if (b[5]) PC = PC+2; //b5
//    if (b[4]) PC = ABUS; //b4
//    if (b[1]) RBUS = AC; //b1
//    if (b[0]) RBUS = ALU_RESULT; //b0
//  end
   
endmodule



